mgc_hls.mgc_io_sync(beh) rtlc_no_parameters
